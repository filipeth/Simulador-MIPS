module mux_jump (endSomador);

endmodule